Simple Resistive Network
v1 0 batt 1.5
r1 batt x 1k
r2 x y 2k
r3 y 0 2k
r4 y 0 3k
.op
.end
